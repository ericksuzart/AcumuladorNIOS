// SistemaEmbarcadoAcumulador_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcadoAcumulador_tb (
	);

	wire         sistemaembarcadoacumulador_inst_clk_bfm_clk_clk;                 // SistemaEmbarcadoAcumulador_inst_clk_bfm:clk -> [SistemaEmbarcadoAcumulador_inst:clk_clk, SistemaEmbarcadoAcumulador_inst_acumulador_conduit_bfm:clk, SistemaEmbarcadoAcumulador_inst_medidordeclock_conduit_bfm:clk, SistemaEmbarcadoAcumulador_inst_reset_bfm:clk]
	wire  [31:0] sistemaembarcadoacumulador_inst_acumulador_conduit_readdata;     // SistemaEmbarcadoAcumulador_inst:acumulador_conduit_readdata -> SistemaEmbarcadoAcumulador_inst_acumulador_conduit_bfm:sig_readdata
	wire  [31:0] sistemaembarcadoacumulador_inst_medidordeclock_conduit_readdata; // SistemaEmbarcadoAcumulador_inst:medidordeclock_conduit_readdata -> SistemaEmbarcadoAcumulador_inst_medidordeclock_conduit_bfm:sig_readdata
	wire         sistemaembarcadoacumulador_inst_reset_bfm_reset_reset;           // SistemaEmbarcadoAcumulador_inst_reset_bfm:reset -> [SistemaEmbarcadoAcumulador_inst:reset_reset_n, SistemaEmbarcadoAcumulador_inst_acumulador_conduit_bfm:reset, SistemaEmbarcadoAcumulador_inst_medidordeclock_conduit_bfm:reset]

	SistemaEmbarcadoAcumulador sistemaembarcadoacumulador_inst (
		.acumulador_conduit_readdata     (sistemaembarcadoacumulador_inst_acumulador_conduit_readdata),     //     acumulador_conduit.readdata
		.clk_clk                         (sistemaembarcadoacumulador_inst_clk_bfm_clk_clk),                 //                    clk.clk
		.medidordeclock_conduit_readdata (sistemaembarcadoacumulador_inst_medidordeclock_conduit_readdata), // medidordeclock_conduit.readdata
		.reset_reset_n                   (sistemaembarcadoacumulador_inst_reset_bfm_reset_reset)            //                  reset.reset_n
	);

	altera_conduit_bfm sistemaembarcadoacumulador_inst_acumulador_conduit_bfm (
		.clk          (sistemaembarcadoacumulador_inst_clk_bfm_clk_clk),             //     clk.clk
		.reset        (~sistemaembarcadoacumulador_inst_reset_bfm_reset_reset),      //   reset.reset
		.sig_readdata (sistemaembarcadoacumulador_inst_acumulador_conduit_readdata)  // conduit.readdata
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sistemaembarcadoacumulador_inst_clk_bfm (
		.clk (sistemaembarcadoacumulador_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm sistemaembarcadoacumulador_inst_medidordeclock_conduit_bfm (
		.clk          (sistemaembarcadoacumulador_inst_clk_bfm_clk_clk),                 //     clk.clk
		.reset        (~sistemaembarcadoacumulador_inst_reset_bfm_reset_reset),          //   reset.reset
		.sig_readdata (sistemaembarcadoacumulador_inst_medidordeclock_conduit_readdata)  // conduit.readdata
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sistemaembarcadoacumulador_inst_reset_bfm (
		.reset (sistemaembarcadoacumulador_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sistemaembarcadoacumulador_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
